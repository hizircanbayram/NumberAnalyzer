library verilog;
use verilog.vl_types.all;
entity numberAnalyzerTestBench is
end numberAnalyzerTestBench;
