library verilog;
use verilog.vl_types.all;
entity isPalindromeTestBench is
end isPalindromeTestBench;
