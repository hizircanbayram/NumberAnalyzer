library verilog;
use verilog.vl_types.all;
entity isFibonacciTestBench is
end isFibonacciTestBench;
