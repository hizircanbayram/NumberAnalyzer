library verilog;
use verilog.vl_types.all;
entity isEvenNumberTestBench is
end isEvenNumberTestBench;
